module mod1

fn init() {}

pub fn say_hi() {
	println('hello from mod1!')
}

pub fn say_hi_str() string {
	return 'hello from mod1!'
}