// E:/Vlang/The_Way_to_V/Chapter_14_V_Modules/owmw module header

module owmw


