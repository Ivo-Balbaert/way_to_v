// E:/Vlang/The_Way_to_V/Chapter_11_Modules_and_Testing/mod1 module header

module mod1


