// sum.v
module sum 

pub fn sum(a, b int) int {
    return a + b
}
