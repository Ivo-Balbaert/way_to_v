module moduleb
 
fn init() {
  println('Initializing module b!')
}

pub fn world() { 
  println('world!') 
} 
