module modulea
 
fn init() {
  println('Initializing module a!')
}

pub fn hello() { 
  print('Hello ') 
} 
